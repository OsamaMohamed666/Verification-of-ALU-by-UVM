`include "seq_item.sv"
`include "base_seq.sv"
`include "direct_seq.sv"
`include "alu_sequencer.sv"
`include "alu_drv.sv"
`include "alu_moni_in.sv"
`include "alu_moni_out.sv"
`include "alu_agent.sv"
`include "alu_sb.sv"
`include "alu_cov.sv"
`include "alu_env.sv"
